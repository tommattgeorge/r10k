import LFSR::*;

typedef LFSR#(t) FeedLFSR#(type t);